module div(
    input wire clk,
    input wire rst,

    input wire [`DataBus] rs1,
    input wire [`DataBus] rs2,

    input wire write_enable,

    output reg [`DataBus] result,
    output reg error 
);

endmodule // div